magic
tech sky130A
timestamp 1636975877
<< nmos >>
rect -99 14 1 514
<< ndiff >>
rect -385 365 -99 514
rect -385 178 -316 365
rect -169 178 -99 365
rect -385 14 -99 178
rect 1 365 287 514
rect 1 178 70 365
rect 217 178 287 365
rect 1 14 287 178
<< ndiffc >>
rect -316 178 -169 365
rect 70 178 217 365
<< poly >>
rect -99 514 1 566
rect -99 -47 1 14
<< locali >>
rect -321 365 -167 400
rect -321 178 -316 365
rect -169 178 -167 365
rect -321 141 -167 178
rect 65 365 219 400
rect 65 178 70 365
rect 217 178 219 365
rect 65 141 219 178
<< end >>
