* SPICE3 file created from (UNNAMED).ext - technology: sky130A

X0 a_1_14# a_n101_n47# a_n385_14# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5.03e+06u l=1.02e+06u
